-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 12.1 Build 243 01/31/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Dec 12 14:42:34 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY JEDA IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        bt : IN STD_LOGIC := '0';
        b1 : IN STD_LOGIC := '0';
        b2 : IN STD_LOGIC := '0';
        b3 : IN STD_LOGIC := '0';
        s1 : IN STD_LOGIC := '0';
        s2 : IN STD_LOGIC := '0';
        s3 : IN STD_LOGIC := '0';
        st : IN STD_LOGIC := '0';
        SM : OUT STD_LOGIC;
        DM : OUT STD_LOGIC
    );
END JEDA;

ARCHITECTURE BEHAVIOR OF JEDA IS
    TYPE type_fstate IS (t,a1,a2,a3,sub1,sub2,sub3,stopup1,stopup2,des1,des2,des3,stopdown1,stopdown2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,bt,b1,b2,b3,s1,s2,s3,st)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= t;
            SM <= '0';
            DM <= '0';
        ELSE
            SM <= '0';
            DM <= '0';
            CASE fstate IS
                WHEN t =>
                    IF ((((NOT((b1 = '1')) AND NOT((b2 = '1'))) AND NOT((b3 = '1'))) AND (bt = '1'))) THEN
                        reg_fstate <= t;
                    ELSIF ((((b1 = '1') AND NOT((bt = '1'))) AND ((b2 = '1') OR (b3 = '1')))) THEN
                        reg_fstate <= sub1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= t;
                    END IF;
                WHEN a1 =>
                    IF (((((b2 = '1') OR (b3 = '1')) AND NOT((b1 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= stopup1;
                    ELSIF (((((b1 = '1') AND NOT((b2 = '1'))) AND NOT((b3 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= a1;
                    ELSIF ((((NOT((b1 = '1')) AND NOT((b2 = '1'))) AND NOT((b3 = '1'))) AND (bt = '1'))) THEN
                        reg_fstate <= stopdown1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= a1;
                    END IF;
                WHEN a2 =>
                    IF (((((b3 = '1') AND NOT((b2 = '1'))) AND NOT((bt = '1'))) AND NOT((b1 = '1')))) THEN
                        reg_fstate <= stopup2;
                    ELSIF ((((NOT((b1 = '1')) AND (b2 = '1')) AND NOT((b3 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= a2;
                    ELSIF (((((b1 = '1') OR (bt = '1')) AND NOT((b2 = '1'))) AND NOT((b3 = '1')))) THEN
                        reg_fstate <= stopdown2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= a2;
                    END IF;
                WHEN a3 =>
                    IF ((((b2 = '1') OR (b1 = '1')) OR (bt = '1'))) THEN
                        reg_fstate <= des3;
                    ELSIF (((((b3 = '1') AND NOT((b1 = '1'))) AND NOT((b2 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= a3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= a3;
                    END IF;
                WHEN sub1 =>
                    IF (((((b1 = '1') AND NOT((b2 = '1'))) AND NOT((b3 = '1'))) AND (s1 = '1'))) THEN
                        reg_fstate <= stopup1;
                    ELSIF ((NOT((b1 = '1')) AND ((b2 = '1') OR (b3 = '1')))) THEN
                        reg_fstate <= sub2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= sub1;
                    END IF;

                    SM <= '1';
                WHEN sub2 =>
                    IF ((((b2 = '1') AND NOT((b3 = '1'))) AND (s2 = '1'))) THEN
                        reg_fstate <= stopup2;
                    ELSIF ((b3 = '1')) THEN
                        reg_fstate <= sub3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= sub2;
                    END IF;

                    SM <= '1';
                WHEN sub3 =>
                    IF (((b3 = '1') AND (s3 = '1'))) THEN
                        reg_fstate <= a3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= sub3;
                    END IF;

                    SM <= '1';
                WHEN stopup1 =>
                    IF (((NOT((b1 = '1')) AND ((b2 = '1') OR (b3 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= sub2;
                    ELSIF (((((b1 = '1') AND NOT((b2 = '1'))) AND NOT((b3 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= a1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= stopup1;
                    END IF;
                WHEN stopup2 =>
                    IF (((((b2 = '1') AND NOT((b3 = '1'))) AND NOT((b1 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= a2;
                    ELSIF ((((NOT((b1 = '1')) AND NOT((b2 = '1'))) AND (b3 = '1')) AND NOT((bt = '1')))) THEN
                        reg_fstate <= sub3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= stopup2;
                    END IF;
                WHEN des1 =>
                    IF ((bt = '1')) THEN
                        reg_fstate <= t;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= des1;
                    END IF;

                    DM <= '1';
                WHEN des2 =>
                    IF ((((((b1 = '1') AND (s1 = '1')) AND NOT((b2 = '1'))) AND NOT((b3 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= stopdown1;
                    ELSIF ((bt = '1')) THEN
                        reg_fstate <= des1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= des2;
                    END IF;

                    DM <= '1';
                WHEN des3 =>
                    IF ((((((b2 = '1') AND (s2 = '1')) AND NOT((b1 = '1'))) AND NOT((b3 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= stopdown2;
                    ELSIF (((b1 = '1') OR (bt = '1'))) THEN
                        reg_fstate <= des2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= des3;
                    END IF;

                    DM <= '1';
                WHEN stopdown1 =>
                    IF (((((b1 = '1') AND NOT((b2 = '1'))) AND NOT((b3 = '1'))) AND NOT((bt = '1')))) THEN
                        reg_fstate <= a1;
                    ELSIF (((bt = '1') AND (st = '1'))) THEN
                        reg_fstate <= des1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= stopdown1;
                    END IF;
                WHEN stopdown2 =>
                    IF (((b1 = '1') OR (bt = '1'))) THEN
                        reg_fstate <= des2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= stopdown2;
                    END IF;
                WHEN OTHERS => 
                    SM <= 'X';
                    DM <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
